LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ADD1 IS 
PORT (
        PCIN: IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
        PCOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
        --QB:OUT STD_LOGIC);
END ADD1;

ARCHITECTURE behav OF ADD1 IS
BEGIN 

	PCout<=PCin+"00000001";
	
  
 
END behav;
