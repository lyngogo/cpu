LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ID IS 
PORT (CLK:IN STD_LOGIC;
        DATAIN: IN  STD_LOGIC;
        DATAOUT:OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
        --QB:OUT STD_LOGIC);
END ID;

ARCHITECTURE behav OF ID IS
BEGIN 

PROCESS (CLK)
    VARIABLE REG8:STD_LOGIC_VECTOR (1 DOWNTO 0);
	  VARIABLE flag:STD_LOGIC ;
BEGIN 
    IF CLK'EVENT AND CLK='1' 
    THEN
        IF flag='0' THEN
              
				REG8(0):=DATAIN;
				flag:='1';
				ELSE   REG8(1):=REG8(0);
				REG8(0):=DATAIN;
				DATAOUT<=REG8;flag:='0'; END IF;
    END IF; 
   
END PROCESS;
END behav;
