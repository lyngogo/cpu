LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY PC IS 
PORT (CLK:IN STD_LOGIC;
        PCIN: IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
        PCOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
        --QB:OUT STD_LOGIC);
END PC;

ARCHITECTURE behav OF PC IS
BEGIN 
PROCESS (CLK)
    VARIABLE REG8:STD_LOGIC_VECTOR (1 DOWNTO 0);
	  VARIABLE flag:STD_LOGIC ;
BEGIN 
    IF CLK'EVENT AND CLK='1' then
		PCOUT<=PCIN;
    END IF; 
   
END PROCESS;
END behav;
